module wand_example(
  input wire a,
  input wire b,
  output wand out
);

  assign out = a;
  assign out = b;

endmodule